module instmem (a,inst);
    input  [31:0] a;
    output [31:0] inst;
    wire   [31:0] rom [0:7];
    assign rom[3'h0] = 32'b00100000000100000000000000010000; // addi  $16, $00, 16    
    assign rom[3'h1] = 32'b00010010000000000000000000000010; // beq   $16, $00, 2     
    assign rom[3'h2] = 32'b00100010000100001111111111111111; // addi  $16, $16, -1    
    assign rom[3'h3] = 32'b00001000000000000000000000000001; // j     0x0001          
    assign rom[3'h4] = 32'b00000000000000000000000000000000; // nop                   
    assign rom[3'h5] = 32'b00000000000000000000000000000000; // nop                   
    assign rom[3'h6] = 32'b00000000000000000000000000000000; // nop                   
    assign rom[3'h7] = 32'b00000000000000000000000000000000; // nop                   
    assign inst = rom[a[4:2]];
endmodule
