//test bench for booth algorithm
module booth4_tb;

//registers for inputs because they hold values
reg [7:0] a, b;
wire [15:0] prod;

//display operands a, b, and product
initial
$monitor ("a = %b, b = %b, prod = %h", a, b, prod);

//apply input vectors
initial
begin
//for examples 6.6 through 6.10
		#0		a = 8'b0001_1011;
				b = 8'b0111_1000;

		#10	a = 8'b1010_1101;
				b = 8'b0011_1110;


		#10	a = 8'b0100_1010;
				b = 8'b1101_1100;

		#10	a = 8'b1010_0010;
				b = 8'b1101_1100;

		#10	a = 8'b0100_1110;
				b = 8'b0010_1011;

//test b[1:0] ---------------------------------------
		#10	a = 8'b1100_1100;
				b = 8'b1100_1100;

		#10	a = 8'b1100_1100;
				b = 8'b1100_1101;

		#10	a = 8'b1100_1100;
				b = 8'b1100_1110;

		#10	a = 8'b1100_1100;
				b = 8'b1100_1111;


//test b[2:1] ---------------------------------------

		#10	a = 8'b0111_1111;
				b = 8'b1011_1000;

		#10	a = 8'b1011_0011;
				b = 8'b1100_1011;

		#10	a = 8'b0111_0000;
				b = 8'b0111_0100;

		#10	a = 8'b0111_0000;
				b = 8'b0111_0110;


//test b[3:2] ---------------------------------------
		#10	a = 8'b0111_1111;
				b = 8'b1011_0000;

		#10	a = 8'b1011_0011;
				b = 8'b1100_0111;

		#10	a = 8'b0111_0000;
				b = 8'b0111_1000;

		#10	a = 8'b0111_0000;
				b = 8'b0111_1110;

//test b[4:3] ---------------------------------------
		#10	a = 8'b0111_1111;
				b = 8'b1010_0000;

		#10	a = 8'b1011_0011;
				b = 8'b1100_1111;

		#10	a = 8'b0111_0000;
				b = 8'b0111_0000;

		#10	a = 8'b0111_0000;
				b = 8'b0111_1110;


//test b[5:4] ---------------------------------------
		#10	a = 8'b0111_1111;
				b = 8'b1000_0000;

		#10	a = 8'b1011_0011;
				b = 8'b1101_1111;

		#10	a = 8'b0111_0000;
				b = 8'b0110_0000;

		#10	a = 8'b0111_0000;
				b = 8'b0111_1110;


//test b[6:5] ---------------------------------------
		#10	a = 8'b0111_1111;
				b = 8'b1000_0000;

		#10	a = 8'b1011_0011;
				b = 8'b1010_1111;

		#10	a = 8'b0111_0000;
				b = 8'b0101_0000;

		#10	a = 8'b0111_0000;
				b = 8'b0111_1110;

//test b[7:6] ---------------------------------------
		#10	a = 8'b0111_1111;
				b = 8'b0010_0000;

		#10	a = 8'b1011_0011;
				b = 8'b0100_1111;

		#10	a = 8'b0111_0000;
				b = 8'b1011_0000;

		#10	a = 8'b0111_0000;
				b = 8'b1111_1110;

		#10	$stop;
end

//instantiate the module into the test bench
booth4 inst1 (
		.a(a),
		.b(b),
		.prod(prod)
		);

endmodule
