module array_multiplier_tb;

reg [31:0] a, b;
wire [31:0] y;

array_multiplier #(
	.width(32)
) uut (
	.a(a),
	.b(b),
	.y(y)
); 

initial begin
    // a = 6
    // b = 9
    // prod = 54
    #10
    a = 32'b00000000000000000000000000000110;
    b = 32'b00000000000000000000000000001001;

    // a = 14
    // b = 12
	// prod = 168
	#10
	a = 32'b00000000000000000000000000001110;
	b = 32'b00000000000000000000000000001100;
		
	// a = 10
	// b = 11
	// prod = 110
	#10
	a = 32'b00000000000000000000000000001010;
	b = 32'b00000000000000000000000000001011;

    // a = 15
	// b = 15
	// prod = 225
	#10
	a = 32'b00000000000000000000000000001111;
	b = 32'b00000000000000000000000000001111;
	
	#10
	$finish;
end

endmodule